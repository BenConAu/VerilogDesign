module DemoModule
begin
  input wire[31:0] in1;
  output reg[31:0] out1;
  case initial
  begin
  end
  case StartState
  begin
  end
  case EndState
  begin
  end
end
