module DemoModule
begin
  case initial
  begin
  end
  case StartState
  begin
  end
  case EndState
  begin
  end
end
