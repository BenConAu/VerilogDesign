module DemoModule
begin
