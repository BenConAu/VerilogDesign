`define MCWaiting   0
`define MCReady     1
`define MCError     2
