module DemoModule
begin
  input wire[7:0] in1;
  output reg[7:0] out1;
  case initial
  begin
  end
  case StartState
  begin
  end
  case EndState
  begin
  end
end
